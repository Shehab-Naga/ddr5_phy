`include "base_test.sv"
`include "ddr_sanity_test.sv"
`include "rand_test.sv"
`include "rand_test_corners.sv"
`include "b2b_test.sv"



