`include "base_seq.sv"
`include "reset_seq.sv"
`include "ddr_sanity_seq.sv"
`include "ACT_seq.sv"
`include "RD_seq.sv"
`include "MRW_seq.sv"
`include "MRR_seq.sv"
`include "PREab_seq.sv"
`include "DES_seq.sv"
`include "dram_resp_seq.sv"
`include "rand_seq.sv"
`include "b2b_seq.sv"
`include "ACT_seq_corners.sv"
`include "RD_seq_corners.sv"
`include "rand_seq_corners.sv"
